LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY PSRModifier_p3_tb IS
END PSRModifier_p3_tb;
 
ARCHITECTURE behavior OF PSRModifier_p3_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT PSRModifier_p3
    PORT(
         rst : IN  std_logic;
         aluop : IN  std_logic_vector(5 downto 0);
         crs1 : IN  std_logic_vector(31 downto 0);
         crs2alu : IN  std_logic_vector(31 downto 0);
         salu : IN  std_logic_vector(31 downto 0);
         nzvc : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '0';
   signal aluop : std_logic_vector(5 downto 0) := (others => '0');
   signal crs1 : std_logic_vector(31 downto 0) := (others => '0');
   signal crs2alu : std_logic_vector(31 downto 0) := (others => '0');
   signal salu : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal nzvc : std_logic_vector(3 downto 0);
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: PSRModifier_p3 PORT MAP (
          rst => rst,
          aluop => aluop,
          crs1 => crs1,
          crs2alu => crs2alu,
          salu => salu,
          nzvc => nzvc
        );
 

   -- Stimulus process
   stim_proc: process
   begin		
      rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "00000000000000000000000001111000";
      wait for 100 ns;	
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "000000";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "000000";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '1';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "011000";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "010000";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "011000";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "011000";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "011000";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "010100";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '1';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010100";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010100";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "000100";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "010100";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "010100";
      salu <= "00000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "011100";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "011100";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "10000000000000000000000001111000";
      crs2alu <= "10000000000000000000000001111000"; 
      aluop <= "011100";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
		rst <= '0';
      crs1 <= "00000000000000000000000001111000";
      crs2alu <= "00000000000000000000000001111000"; 
      aluop <= "011100";
      salu <= "10000000000000000000000000000000";
      wait for 100 ns;
   end process;

END;

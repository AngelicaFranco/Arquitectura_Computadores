library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity InstructionMemory_p1 is
    Port ( rst : in  STD_LOGIC;
           pc : in  STD_LOGIC_VECTOR (31 downto 0);
           instructionout : out  STD_LOGIC_VECTOR (31 downto 0));
end InstructionMemory_p1;

architecture Behavioral of InstructionMemory_p1 is
	type rom_type is array (0 to 63) of STD_LOGIC_VECTOR (31 downto 0);
	signal instructions : rom_type := (X"01000000",
												  "00010000100000000000000000001110",
												  X"01000000",
												  "10100000000100000010000000000000",
												  "10100010000100000010000000000000",
												  "10000000101001000100000000011001",
												  "00010110100000000000000000000111",
												  X"01000000",
												  "10100100000001000000000000011000",
												  "10100000000100000000000000010010",
												  "10100100000001000110000000000001",
												  "00010000101111111111111111111010",
												  "10100010000100000000000000010010",
												  "10000001110000111110000000000010", 
												  "10010000000100000000000000010000", 
												  "10110000000100000010000000000011",  -- X
												  "10110010000100000010000000001000", -- Y
												  "01111111111111111111111111110010", 
												  X"01000000", X"01000000",
												  "10010010000100000000000000001000",  
												  X"01000000", X"01000000", X"01000000",  
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000", 
												  X"01000000", X"01000000", X"01000000", X"01000000");
	
begin
	process (rst, pc)
		begin
			if (rst = '1') then
				instructionout <= (others => '0');
			else
				instructionout <= instructions(conv_integer(pc(5 downto 0)));
			end if;
	end process;
end Behavioral;

